`timescale 10 ns / 1 ns