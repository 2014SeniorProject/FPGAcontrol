`define debug