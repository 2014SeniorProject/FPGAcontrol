module MotorControl_TB(

    );